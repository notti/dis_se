library IEEE;
        use IEEE.STD_LOGIC_1164.ALL;
        use IEEE.NUMERIC_STD.ALL;
library std;
        use std.textio.all;

library work;
        use work.all;
        use work.procedures.all;

entity tb_mp is
end tb_mp;


architecture behav of tb_mp is
       signal rst     :  std_logic := '1';
       signal clk     :  std_logic := '0';
       signal pdata   :  t_data2 := (others => '0');
       signal pdata_rd : std_logic := '0';
       signal start   :  std_logic := '0';
       signal busy    :  std_logic := '0';
       signal mem_addra :  std_logic_vector(9 downto 0) := (others => '0'); 
       signal mem_ena   :  std_logic := '0';
       signal mem_doa :  t_data := (others => '0');
       signal mem_addrb :  std_logic_vector(9 downto 0) := (others => '0'); 
       signal mem_enb   :  std_logic := '0';
       signal mem_dob :  t_data := (others => '0');
       signal reg_addra:  t_data := (others => '0');
       signal reg_ena  :  std_logic := '0';
       signal reg_doa  :  t_data := (others => '0');
       signal reg_addrb:  t_data := (others => '0');
       signal reg_enb  :  std_logic := '0';
       signal reg_dob  :  t_data := (others => '0');
       signal clk2x   : std_logic := '0';


       procedure prog_cmd(cmd     : in t_vliw;
                        which     : in natural;
                        signal start   : out std_logic;
                        signal pdata   : out t_data2) is
           variable tmp : std_logic_vector(VLIW_HIGH downto 0);
       begin
           tmp := vliw2slv(cmd);
           start <= '1';
           pdata <= "1111111111111" & std_logic_vector(to_unsigned(which, 3));
           wait for 20 ns;
           start <= '0';
           for i in 0 to VLIW_HIGH/16-1 loop
               pdata <= tmp((i+1)*16-1 downto i*16);
               wait for 20 ns;
           end loop;
           pdata(VLIW_HIGH mod 8 downto 0) <= tmp(VLIW_HIGH downto (VLIW_HIGH/16)*16);
           wait for 40 ns;
       end procedure;

       type int_arr is array(natural range <>) of integer;
       signal sine_wave : int_arr(0 to 255) := (0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0, -26, -52, -75, -95, -110, -121, -127, -127, -121, -110, -95, -75, -52, -26, 0, 26, 52, 75, 95, 110, 121, 127, 127, 121, 110, 95, 75, 52, 26, 0);

       type int_arr_arr is array(natural range <>) of int_arr(0 to 3);
       signal bflys : int_arr_arr(0 to 1023) := (
            (0, 1, 64, 0),
            (2, 3, 64, 0),
            (4, 5, 64, 0),
            (6, 7, 64, 0),
            (8, 9, 64, 0),
            (10, 11, 64, 0),
            (12, 13, 64, 0),
            (14, 15, 64, 0),
            (16, 17, 64, 0),
            (18, 19, 64, 0),
            (20, 21, 64, 0),
            (22, 23, 64, 0),
            (24, 25, 64, 0),
            (26, 27, 64, 0),
            (28, 29, 64, 0),
            (30, 31, 64, 0),
            (32, 33, 64, 0),
            (34, 35, 64, 0),
            (36, 37, 64, 0),
            (38, 39, 64, 0),
            (40, 41, 64, 0),
            (42, 43, 64, 0),
            (44, 45, 64, 0),
            (46, 47, 64, 0),
            (48, 49, 64, 0),
            (50, 51, 64, 0),
            (52, 53, 64, 0),
            (54, 55, 64, 0),
            (56, 57, 64, 0),
            (58, 59, 64, 0),
            (60, 61, 64, 0),
            (62, 63, 64, 0),
            (64, 65, 64, 0),
            (66, 67, 64, 0),
            (68, 69, 64, 0),
            (70, 71, 64, 0),
            (72, 73, 64, 0),
            (74, 75, 64, 0),
            (76, 77, 64, 0),
            (78, 79, 64, 0),
            (80, 81, 64, 0),
            (82, 83, 64, 0),
            (84, 85, 64, 0),
            (86, 87, 64, 0),
            (88, 89, 64, 0),
            (90, 91, 64, 0),
            (92, 93, 64, 0),
            (94, 95, 64, 0),
            (96, 97, 64, 0),
            (98, 99, 64, 0),
            (100, 101, 64, 0),
            (102, 103, 64, 0),
            (104, 105, 64, 0),
            (106, 107, 64, 0),
            (108, 109, 64, 0),
            (110, 111, 64, 0),
            (112, 113, 64, 0),
            (114, 115, 64, 0),
            (116, 117, 64, 0),
            (118, 119, 64, 0),
            (120, 121, 64, 0),
            (122, 123, 64, 0),
            (124, 125, 64, 0),
            (126, 127, 64, 0),
            (128, 129, 64, 0),
            (130, 131, 64, 0),
            (132, 133, 64, 0),
            (134, 135, 64, 0),
            (136, 137, 64, 0),
            (138, 139, 64, 0),
            (140, 141, 64, 0),
            (142, 143, 64, 0),
            (144, 145, 64, 0),
            (146, 147, 64, 0),
            (148, 149, 64, 0),
            (150, 151, 64, 0),
            (152, 153, 64, 0),
            (154, 155, 64, 0),
            (156, 157, 64, 0),
            (158, 159, 64, 0),
            (160, 161, 64, 0),
            (162, 163, 64, 0),
            (164, 165, 64, 0),
            (166, 167, 64, 0),
            (168, 169, 64, 0),
            (170, 171, 64, 0),
            (172, 173, 64, 0),
            (174, 175, 64, 0),
            (176, 177, 64, 0),
            (178, 179, 64, 0),
            (180, 181, 64, 0),
            (182, 183, 64, 0),
            (184, 185, 64, 0),
            (186, 187, 64, 0),
            (188, 189, 64, 0),
            (190, 191, 64, 0),
            (192, 193, 64, 0),
            (194, 195, 64, 0),
            (196, 197, 64, 0),
            (198, 199, 64, 0),
            (200, 201, 64, 0),
            (202, 203, 64, 0),
            (204, 205, 64, 0),
            (206, 207, 64, 0),
            (208, 209, 64, 0),
            (210, 211, 64, 0),
            (212, 213, 64, 0),
            (214, 215, 64, 0),
            (216, 217, 64, 0),
            (218, 219, 64, 0),
            (220, 221, 64, 0),
            (222, 223, 64, 0),
            (224, 225, 64, 0),
            (226, 227, 64, 0),
            (228, 229, 64, 0),
            (230, 231, 64, 0),
            (232, 233, 64, 0),
            (234, 235, 64, 0),
            (236, 237, 64, 0),
            (238, 239, 64, 0),
            (240, 241, 64, 0),
            (242, 243, 64, 0),
            (244, 245, 64, 0),
            (246, 247, 64, 0),
            (248, 249, 64, 0),
            (250, 251, 64, 0),
            (252, 253, 64, 0),
            (254, 255, 64, 0),
            (0, 2, 64, 0),
            (4, 6, 64, 0),
            (8, 10, 64, 0),
            (12, 14, 64, 0),
            (16, 18, 64, 0),
            (20, 22, 64, 0),
            (24, 26, 64, 0),
            (28, 30, 64, 0),
            (32, 34, 64, 0),
            (36, 38, 64, 0),
            (40, 42, 64, 0),
            (44, 46, 64, 0),
            (48, 50, 64, 0),
            (52, 54, 64, 0),
            (56, 58, 64, 0),
            (60, 62, 64, 0),
            (64, 66, 64, 0),
            (68, 70, 64, 0),
            (72, 74, 64, 0),
            (76, 78, 64, 0),
            (80, 82, 64, 0),
            (84, 86, 64, 0),
            (88, 90, 64, 0),
            (92, 94, 64, 0),
            (96, 98, 64, 0),
            (100, 102, 64, 0),
            (104, 106, 64, 0),
            (108, 110, 64, 0),
            (112, 114, 64, 0),
            (116, 118, 64, 0),
            (120, 122, 64, 0),
            (124, 126, 64, 0),
            (128, 130, 64, 0),
            (132, 134, 64, 0),
            (136, 138, 64, 0),
            (140, 142, 64, 0),
            (144, 146, 64, 0),
            (148, 150, 64, 0),
            (152, 154, 64, 0),
            (156, 158, 64, 0),
            (160, 162, 64, 0),
            (164, 166, 64, 0),
            (168, 170, 64, 0),
            (172, 174, 64, 0),
            (176, 178, 64, 0),
            (180, 182, 64, 0),
            (184, 186, 64, 0),
            (188, 190, 64, 0),
            (192, 194, 64, 0),
            (196, 198, 64, 0),
            (200, 202, 64, 0),
            (204, 206, 64, 0),
            (208, 210, 64, 0),
            (212, 214, 64, 0),
            (216, 218, 64, 0),
            (220, 222, 64, 0),
            (224, 226, 64, 0),
            (228, 230, 64, 0),
            (232, 234, 64, 0),
            (236, 238, 64, 0),
            (240, 242, 64, 0),
            (244, 246, 64, 0),
            (248, 250, 64, 0),
            (252, 254, 64, 0),
            (1, 3, 0, -64),
            (5, 7, 0, -64),
            (9, 11, 0, -64),
            (13, 15, 0, -64),
            (17, 19, 0, -64),
            (21, 23, 0, -64),
            (25, 27, 0, -64),
            (29, 31, 0, -64),
            (33, 35, 0, -64),
            (37, 39, 0, -64),
            (41, 43, 0, -64),
            (45, 47, 0, -64),
            (49, 51, 0, -64),
            (53, 55, 0, -64),
            (57, 59, 0, -64),
            (61, 63, 0, -64),
            (65, 67, 0, -64),
            (69, 71, 0, -64),
            (73, 75, 0, -64),
            (77, 79, 0, -64),
            (81, 83, 0, -64),
            (85, 87, 0, -64),
            (89, 91, 0, -64),
            (93, 95, 0, -64),
            (97, 99, 0, -64),
            (101, 103, 0, -64),
            (105, 107, 0, -64),
            (109, 111, 0, -64),
            (113, 115, 0, -64),
            (117, 119, 0, -64),
            (121, 123, 0, -64),
            (125, 127, 0, -64),
            (129, 131, 0, -64),
            (133, 135, 0, -64),
            (137, 139, 0, -64),
            (141, 143, 0, -64),
            (145, 147, 0, -64),
            (149, 151, 0, -64),
            (153, 155, 0, -64),
            (157, 159, 0, -64),
            (161, 163, 0, -64),
            (165, 167, 0, -64),
            (169, 171, 0, -64),
            (173, 175, 0, -64),
            (177, 179, 0, -64),
            (181, 183, 0, -64),
            (185, 187, 0, -64),
            (189, 191, 0, -64),
            (193, 195, 0, -64),
            (197, 199, 0, -64),
            (201, 203, 0, -64),
            (205, 207, 0, -64),
            (209, 211, 0, -64),
            (213, 215, 0, -64),
            (217, 219, 0, -64),
            (221, 223, 0, -64),
            (225, 227, 0, -64),
            (229, 231, 0, -64),
            (233, 235, 0, -64),
            (237, 239, 0, -64),
            (241, 243, 0, -64),
            (245, 247, 0, -64),
            (249, 251, 0, -64),
            (253, 255, 0, -64),
            (0, 4, 64, 0),
            (8, 12, 64, 0),
            (16, 20, 64, 0),
            (24, 28, 64, 0),
            (32, 36, 64, 0),
            (40, 44, 64, 0),
            (48, 52, 64, 0),
            (56, 60, 64, 0),
            (64, 68, 64, 0),
            (72, 76, 64, 0),
            (80, 84, 64, 0),
            (88, 92, 64, 0),
            (96, 100, 64, 0),
            (104, 108, 64, 0),
            (112, 116, 64, 0),
            (120, 124, 64, 0),
            (128, 132, 64, 0),
            (136, 140, 64, 0),
            (144, 148, 64, 0),
            (152, 156, 64, 0),
            (160, 164, 64, 0),
            (168, 172, 64, 0),
            (176, 180, 64, 0),
            (184, 188, 64, 0),
            (192, 196, 64, 0),
            (200, 204, 64, 0),
            (208, 212, 64, 0),
            (216, 220, 64, 0),
            (224, 228, 64, 0),
            (232, 236, 64, 0),
            (240, 244, 64, 0),
            (248, 252, 64, 0),
            (1, 5, 45, -45),
            (9, 13, 45, -45),
            (17, 21, 45, -45),
            (25, 29, 45, -45),
            (33, 37, 45, -45),
            (41, 45, 45, -45),
            (49, 53, 45, -45),
            (57, 61, 45, -45),
            (65, 69, 45, -45),
            (73, 77, 45, -45),
            (81, 85, 45, -45),
            (89, 93, 45, -45),
            (97, 101, 45, -45),
            (105, 109, 45, -45),
            (113, 117, 45, -45),
            (121, 125, 45, -45),
            (129, 133, 45, -45),
            (137, 141, 45, -45),
            (145, 149, 45, -45),
            (153, 157, 45, -45),
            (161, 165, 45, -45),
            (169, 173, 45, -45),
            (177, 181, 45, -45),
            (185, 189, 45, -45),
            (193, 197, 45, -45),
            (201, 205, 45, -45),
            (209, 213, 45, -45),
            (217, 221, 45, -45),
            (225, 229, 45, -45),
            (233, 237, 45, -45),
            (241, 245, 45, -45),
            (249, 253, 45, -45),
            (2, 6, 0, -64),
            (10, 14, 0, -64),
            (18, 22, 0, -64),
            (26, 30, 0, -64),
            (34, 38, 0, -64),
            (42, 46, 0, -64),
            (50, 54, 0, -64),
            (58, 62, 0, -64),
            (66, 70, 0, -64),
            (74, 78, 0, -64),
            (82, 86, 0, -64),
            (90, 94, 0, -64),
            (98, 102, 0, -64),
            (106, 110, 0, -64),
            (114, 118, 0, -64),
            (122, 126, 0, -64),
            (130, 134, 0, -64),
            (138, 142, 0, -64),
            (146, 150, 0, -64),
            (154, 158, 0, -64),
            (162, 166, 0, -64),
            (170, 174, 0, -64),
            (178, 182, 0, -64),
            (186, 190, 0, -64),
            (194, 198, 0, -64),
            (202, 206, 0, -64),
            (210, 214, 0, -64),
            (218, 222, 0, -64),
            (226, 230, 0, -64),
            (234, 238, 0, -64),
            (242, 246, 0, -64),
            (250, 254, 0, -64),
            (3, 7, -45, -45),
            (11, 15, -45, -45),
            (19, 23, -45, -45),
            (27, 31, -45, -45),
            (35, 39, -45, -45),
            (43, 47, -45, -45),
            (51, 55, -45, -45),
            (59, 63, -45, -45),
            (67, 71, -45, -45),
            (75, 79, -45, -45),
            (83, 87, -45, -45),
            (91, 95, -45, -45),
            (99, 103, -45, -45),
            (107, 111, -45, -45),
            (115, 119, -45, -45),
            (123, 127, -45, -45),
            (131, 135, -45, -45),
            (139, 143, -45, -45),
            (147, 151, -45, -45),
            (155, 159, -45, -45),
            (163, 167, -45, -45),
            (171, 175, -45, -45),
            (179, 183, -45, -45),
            (187, 191, -45, -45),
            (195, 199, -45, -45),
            (203, 207, -45, -45),
            (211, 215, -45, -45),
            (219, 223, -45, -45),
            (227, 231, -45, -45),
            (235, 239, -45, -45),
            (243, 247, -45, -45),
            (251, 255, -45, -45),
            (0, 8, 64, 0),
            (16, 24, 64, 0),
            (32, 40, 64, 0),
            (48, 56, 64, 0),
            (64, 72, 64, 0),
            (80, 88, 64, 0),
            (96, 104, 64, 0),
            (112, 120, 64, 0),
            (128, 136, 64, 0),
            (144, 152, 64, 0),
            (160, 168, 64, 0),
            (176, 184, 64, 0),
            (192, 200, 64, 0),
            (208, 216, 64, 0),
            (224, 232, 64, 0),
            (240, 248, 64, 0),
            (1, 9, 59, -24),
            (17, 25, 59, -24),
            (33, 41, 59, -24),
            (49, 57, 59, -24),
            (65, 73, 59, -24),
            (81, 89, 59, -24),
            (97, 105, 59, -24),
            (113, 121, 59, -24),
            (129, 137, 59, -24),
            (145, 153, 59, -24),
            (161, 169, 59, -24),
            (177, 185, 59, -24),
            (193, 201, 59, -24),
            (209, 217, 59, -24),
            (225, 233, 59, -24),
            (241, 249, 59, -24),
            (2, 10, 45, -45),
            (18, 26, 45, -45),
            (34, 42, 45, -45),
            (50, 58, 45, -45),
            (66, 74, 45, -45),
            (82, 90, 45, -45),
            (98, 106, 45, -45),
            (114, 122, 45, -45),
            (130, 138, 45, -45),
            (146, 154, 45, -45),
            (162, 170, 45, -45),
            (178, 186, 45, -45),
            (194, 202, 45, -45),
            (210, 218, 45, -45),
            (226, 234, 45, -45),
            (242, 250, 45, -45),
            (3, 11, 24, -59),
            (19, 27, 24, -59),
            (35, 43, 24, -59),
            (51, 59, 24, -59),
            (67, 75, 24, -59),
            (83, 91, 24, -59),
            (99, 107, 24, -59),
            (115, 123, 24, -59),
            (131, 139, 24, -59),
            (147, 155, 24, -59),
            (163, 171, 24, -59),
            (179, 187, 24, -59),
            (195, 203, 24, -59),
            (211, 219, 24, -59),
            (227, 235, 24, -59),
            (243, 251, 24, -59),
            (4, 12, 0, -64),
            (20, 28, 0, -64),
            (36, 44, 0, -64),
            (52, 60, 0, -64),
            (68, 76, 0, -64),
            (84, 92, 0, -64),
            (100, 108, 0, -64),
            (116, 124, 0, -64),
            (132, 140, 0, -64),
            (148, 156, 0, -64),
            (164, 172, 0, -64),
            (180, 188, 0, -64),
            (196, 204, 0, -64),
            (212, 220, 0, -64),
            (228, 236, 0, -64),
            (244, 252, 0, -64),
            (5, 13, -24, -59),
            (21, 29, -24, -59),
            (37, 45, -24, -59),
            (53, 61, -24, -59),
            (69, 77, -24, -59),
            (85, 93, -24, -59),
            (101, 109, -24, -59),
            (117, 125, -24, -59),
            (133, 141, -24, -59),
            (149, 157, -24, -59),
            (165, 173, -24, -59),
            (181, 189, -24, -59),
            (197, 205, -24, -59),
            (213, 221, -24, -59),
            (229, 237, -24, -59),
            (245, 253, -24, -59),
            (6, 14, -45, -45),
            (22, 30, -45, -45),
            (38, 46, -45, -45),
            (54, 62, -45, -45),
            (70, 78, -45, -45),
            (86, 94, -45, -45),
            (102, 110, -45, -45),
            (118, 126, -45, -45),
            (134, 142, -45, -45),
            (150, 158, -45, -45),
            (166, 174, -45, -45),
            (182, 190, -45, -45),
            (198, 206, -45, -45),
            (214, 222, -45, -45),
            (230, 238, -45, -45),
            (246, 254, -45, -45),
            (7, 15, -59, -24),
            (23, 31, -59, -24),
            (39, 47, -59, -24),
            (55, 63, -59, -24),
            (71, 79, -59, -24),
            (87, 95, -59, -24),
            (103, 111, -59, -24),
            (119, 127, -59, -24),
            (135, 143, -59, -24),
            (151, 159, -59, -24),
            (167, 175, -59, -24),
            (183, 191, -59, -24),
            (199, 207, -59, -24),
            (215, 223, -59, -24),
            (231, 239, -59, -24),
            (247, 255, -59, -24),
            (0, 16, 64, 0),
            (32, 48, 64, 0),
            (64, 80, 64, 0),
            (96, 112, 64, 0),
            (128, 144, 64, 0),
            (160, 176, 64, 0),
            (192, 208, 64, 0),
            (224, 240, 64, 0),
            (1, 17, 62, -12),
            (33, 49, 62, -12),
            (65, 81, 62, -12),
            (97, 113, 62, -12),
            (129, 145, 62, -12),
            (161, 177, 62, -12),
            (193, 209, 62, -12),
            (225, 241, 62, -12),
            (2, 18, 59, -24),
            (34, 50, 59, -24),
            (66, 82, 59, -24),
            (98, 114, 59, -24),
            (130, 146, 59, -24),
            (162, 178, 59, -24),
            (194, 210, 59, -24),
            (226, 242, 59, -24),
            (3, 19, 53, -36),
            (35, 51, 53, -36),
            (67, 83, 53, -36),
            (99, 115, 53, -36),
            (131, 147, 53, -36),
            (163, 179, 53, -36),
            (195, 211, 53, -36),
            (227, 243, 53, -36),
            (4, 20, 45, -45),
            (36, 52, 45, -45),
            (68, 84, 45, -45),
            (100, 116, 45, -45),
            (132, 148, 45, -45),
            (164, 180, 45, -45),
            (196, 212, 45, -45),
            (228, 244, 45, -45),
            (5, 21, 35, -53),
            (37, 53, 35, -53),
            (69, 85, 35, -53),
            (101, 117, 35, -53),
            (133, 149, 35, -53),
            (165, 181, 35, -53),
            (197, 213, 35, -53),
            (229, 245, 35, -53),
            (6, 22, 24, -59),
            (38, 54, 24, -59),
            (70, 86, 24, -59),
            (102, 118, 24, -59),
            (134, 150, 24, -59),
            (166, 182, 24, -59),
            (198, 214, 24, -59),
            (230, 246, 24, -59),
            (7, 23, 12, -63),
            (39, 55, 12, -63),
            (71, 87, 12, -63),
            (103, 119, 12, -63),
            (135, 151, 12, -63),
            (167, 183, 12, -63),
            (199, 215, 12, -63),
            (231, 247, 12, -63),
            (8, 24, 0, -64),
            (40, 56, 0, -64),
            (72, 88, 0, -64),
            (104, 120, 0, -64),
            (136, 152, 0, -64),
            (168, 184, 0, -64),
            (200, 216, 0, -64),
            (232, 248, 0, -64),
            (9, 25, -12, -63),
            (41, 57, -12, -63),
            (73, 89, -12, -63),
            (105, 121, -12, -63),
            (137, 153, -12, -63),
            (169, 185, -12, -63),
            (201, 217, -12, -63),
            (233, 249, -12, -63),
            (10, 26, -24, -59),
            (42, 58, -24, -59),
            (74, 90, -24, -59),
            (106, 122, -24, -59),
            (138, 154, -24, -59),
            (170, 186, -24, -59),
            (202, 218, -24, -59),
            (234, 250, -24, -59),
            (11, 27, -36, -53),
            (43, 59, -36, -53),
            (75, 91, -36, -53),
            (107, 123, -36, -53),
            (139, 155, -36, -53),
            (171, 187, -36, -53),
            (203, 219, -36, -53),
            (235, 251, -36, -53),
            (12, 28, -45, -45),
            (44, 60, -45, -45),
            (76, 92, -45, -45),
            (108, 124, -45, -45),
            (140, 156, -45, -45),
            (172, 188, -45, -45),
            (204, 220, -45, -45),
            (236, 252, -45, -45),
            (13, 29, -53, -36),
            (45, 61, -53, -36),
            (77, 93, -53, -36),
            (109, 125, -53, -36),
            (141, 157, -53, -36),
            (173, 189, -53, -36),
            (205, 221, -53, -36),
            (237, 253, -53, -36),
            (14, 30, -59, -24),
            (46, 62, -59, -24),
            (78, 94, -59, -24),
            (110, 126, -59, -24),
            (142, 158, -59, -24),
            (174, 190, -59, -24),
            (206, 222, -59, -24),
            (238, 254, -59, -24),
            (15, 31, -63, -12),
            (47, 63, -63, -12),
            (79, 95, -63, -12),
            (111, 127, -63, -12),
            (143, 159, -63, -12),
            (175, 191, -63, -12),
            (207, 223, -63, -12),
            (239, 255, -63, -12),
            (0, 32, 64, 0),
            (64, 96, 64, 0),
            (128, 160, 64, 0),
            (192, 224, 64, 0),
            (1, 33, 63, -6),
            (65, 97, 63, -6),
            (129, 161, 63, -6),
            (193, 225, 63, -6),
            (2, 34, 62, -12),
            (66, 98, 62, -12),
            (130, 162, 62, -12),
            (194, 226, 62, -12),
            (3, 35, 61, -19),
            (67, 99, 61, -19),
            (131, 163, 61, -19),
            (195, 227, 61, -19),
            (4, 36, 59, -24),
            (68, 100, 59, -24),
            (132, 164, 59, -24),
            (196, 228, 59, -24),
            (5, 37, 56, -30),
            (69, 101, 56, -30),
            (133, 165, 56, -30),
            (197, 229, 56, -30),
            (6, 38, 53, -36),
            (70, 102, 53, -36),
            (134, 166, 53, -36),
            (198, 230, 53, -36),
            (7, 39, 49, -41),
            (71, 103, 49, -41),
            (135, 167, 49, -41),
            (199, 231, 49, -41),
            (8, 40, 45, -45),
            (72, 104, 45, -45),
            (136, 168, 45, -45),
            (200, 232, 45, -45),
            (9, 41, 40, -49),
            (73, 105, 40, -49),
            (137, 169, 40, -49),
            (201, 233, 40, -49),
            (10, 42, 35, -53),
            (74, 106, 35, -53),
            (138, 170, 35, -53),
            (202, 234, 35, -53),
            (11, 43, 30, -56),
            (75, 107, 30, -56),
            (139, 171, 30, -56),
            (203, 235, 30, -56),
            (12, 44, 24, -59),
            (76, 108, 24, -59),
            (140, 172, 24, -59),
            (204, 236, 24, -59),
            (13, 45, 18, -61),
            (77, 109, 18, -61),
            (141, 173, 18, -61),
            (205, 237, 18, -61),
            (14, 46, 12, -63),
            (78, 110, 12, -63),
            (142, 174, 12, -63),
            (206, 238, 12, -63),
            (15, 47, 6, -64),
            (79, 111, 6, -64),
            (143, 175, 6, -64),
            (207, 239, 6, -64),
            (16, 48, 0, -64),
            (80, 112, 0, -64),
            (144, 176, 0, -64),
            (208, 240, 0, -64),
            (17, 49, -6, -64),
            (81, 113, -6, -64),
            (145, 177, -6, -64),
            (209, 241, -6, -64),
            (18, 50, -12, -63),
            (82, 114, -12, -63),
            (146, 178, -12, -63),
            (210, 242, -12, -63),
            (19, 51, -19, -61),
            (83, 115, -19, -61),
            (147, 179, -19, -61),
            (211, 243, -19, -61),
            (20, 52, -24, -59),
            (84, 116, -24, -59),
            (148, 180, -24, -59),
            (212, 244, -24, -59),
            (21, 53, -30, -56),
            (85, 117, -30, -56),
            (149, 181, -30, -56),
            (213, 245, -30, -56),
            (22, 54, -36, -53),
            (86, 118, -36, -53),
            (150, 182, -36, -53),
            (214, 246, -36, -53),
            (23, 55, -41, -49),
            (87, 119, -41, -49),
            (151, 183, -41, -49),
            (215, 247, -41, -49),
            (24, 56, -45, -45),
            (88, 120, -45, -45),
            (152, 184, -45, -45),
            (216, 248, -45, -45),
            (25, 57, -49, -41),
            (89, 121, -49, -41),
            (153, 185, -49, -41),
            (217, 249, -49, -41),
            (26, 58, -53, -36),
            (90, 122, -53, -36),
            (154, 186, -53, -36),
            (218, 250, -53, -36),
            (27, 59, -56, -30),
            (91, 123, -56, -30),
            (155, 187, -56, -30),
            (219, 251, -56, -30),
            (28, 60, -59, -24),
            (92, 124, -59, -24),
            (156, 188, -59, -24),
            (220, 252, -59, -24),
            (29, 61, -61, -19),
            (93, 125, -61, -19),
            (157, 189, -61, -19),
            (221, 253, -61, -19),
            (30, 62, -63, -12),
            (94, 126, -63, -12),
            (158, 190, -63, -12),
            (222, 254, -63, -12),
            (31, 63, -64, -6),
            (95, 127, -64, -6),
            (159, 191, -64, -6),
            (223, 255, -64, -6),
            (0, 64, 64, 0),
            (128, 192, 64, 0),
            (1, 65, 63, -3),
            (129, 193, 63, -3),
            (2, 66, 63, -6),
            (130, 194, 63, -6),
            (3, 67, 63, -9),
            (131, 195, 63, -9),
            (4, 68, 62, -12),
            (132, 196, 62, -12),
            (5, 69, 62, -16),
            (133, 197, 62, -16),
            (6, 70, 61, -19),
            (134, 198, 61, -19),
            (7, 71, 60, -22),
            (135, 199, 60, -22),
            (8, 72, 59, -24),
            (136, 200, 59, -24),
            (9, 73, 57, -27),
            (137, 201, 57, -27),
            (10, 74, 56, -30),
            (138, 202, 56, -30),
            (11, 75, 54, -33),
            (139, 203, 54, -33),
            (12, 76, 53, -36),
            (140, 204, 53, -36),
            (13, 77, 51, -38),
            (141, 205, 51, -38),
            (14, 78, 49, -41),
            (142, 206, 49, -41),
            (15, 79, 47, -43),
            (143, 207, 47, -43),
            (16, 80, 45, -45),
            (144, 208, 45, -45),
            (17, 81, 42, -47),
            (145, 209, 42, -47),
            (18, 82, 40, -49),
            (146, 210, 40, -49),
            (19, 83, 38, -51),
            (147, 211, 38, -51),
            (20, 84, 35, -53),
            (148, 212, 35, -53),
            (21, 85, 32, -55),
            (149, 213, 32, -55),
            (22, 86, 30, -56),
            (150, 214, 30, -56),
            (23, 87, 27, -58),
            (151, 215, 27, -58),
            (24, 88, 24, -59),
            (152, 216, 24, -59),
            (25, 89, 21, -60),
            (153, 217, 21, -60),
            (26, 90, 18, -61),
            (154, 218, 18, -61),
            (27, 91, 15, -62),
            (155, 219, 15, -62),
            (28, 92, 12, -63),
            (156, 220, 12, -63),
            (29, 93, 9, -63),
            (157, 221, 9, -63),
            (30, 94, 6, -64),
            (158, 222, 6, -64),
            (31, 95, 3, -64),
            (159, 223, 3, -64),
            (32, 96, 0, -64),
            (160, 224, 0, -64),
            (33, 97, -3, -64),
            (161, 225, -3, -64),
            (34, 98, -6, -64),
            (162, 226, -6, -64),
            (35, 99, -9, -63),
            (163, 227, -9, -63),
            (36, 100, -12, -63),
            (164, 228, -12, -63),
            (37, 101, -16, -62),
            (165, 229, -16, -62),
            (38, 102, -19, -61),
            (166, 230, -19, -61),
            (39, 103, -22, -60),
            (167, 231, -22, -60),
            (40, 104, -24, -59),
            (168, 232, -24, -59),
            (41, 105, -27, -58),
            (169, 233, -27, -58),
            (42, 106, -30, -56),
            (170, 234, -30, -56),
            (43, 107, -33, -55),
            (171, 235, -33, -55),
            (44, 108, -36, -53),
            (172, 236, -36, -53),
            (45, 109, -38, -51),
            (173, 237, -38, -51),
            (46, 110, -41, -49),
            (174, 238, -41, -49),
            (47, 111, -43, -47),
            (175, 239, -43, -47),
            (48, 112, -45, -45),
            (176, 240, -45, -45),
            (49, 113, -47, -43),
            (177, 241, -47, -43),
            (50, 114, -49, -41),
            (178, 242, -49, -41),
            (51, 115, -51, -38),
            (179, 243, -51, -38),
            (52, 116, -53, -36),
            (180, 244, -53, -36),
            (53, 117, -55, -33),
            (181, 245, -55, -33),
            (54, 118, -56, -30),
            (182, 246, -56, -30),
            (55, 119, -58, -27),
            (183, 247, -58, -27),
            (56, 120, -59, -24),
            (184, 248, -59, -24),
            (57, 121, -60, -22),
            (185, 249, -60, -22),
            (58, 122, -61, -19),
            (186, 250, -61, -19),
            (59, 123, -62, -16),
            (187, 251, -62, -16),
            (60, 124, -63, -12),
            (188, 252, -63, -12),
            (61, 125, -63, -9),
            (189, 253, -63, -9),
            (62, 126, -64, -6),
            (190, 254, -64, -6),
            (63, 127, -64, -3),
            (191, 255, -64, -3),
            (0, 128, 64, 0),
            (1, 129, 63, -2),
            (2, 130, 63, -3),
            (3, 131, 63, -5),
            (4, 132, 63, -6),
            (5, 133, 63, -8),
            (6, 134, 63, -9),
            (7, 135, 63, -11),
            (8, 136, 62, -12),
            (9, 137, 62, -14),
            (10, 138, 62, -16),
            (11, 139, 61, -17),
            (12, 140, 61, -19),
            (13, 141, 60, -20),
            (14, 142, 60, -22),
            (15, 143, 59, -23),
            (16, 144, 59, -24),
            (17, 145, 58, -26),
            (18, 146, 57, -27),
            (19, 147, 57, -29),
            (20, 148, 56, -30),
            (21, 149, 55, -32),
            (22, 150, 54, -33),
            (23, 151, 54, -34),
            (24, 152, 53, -36),
            (25, 153, 52, -37),
            (26, 154, 51, -38),
            (27, 155, 50, -39),
            (28, 156, 49, -41),
            (29, 157, 48, -42),
            (30, 158, 47, -43),
            (31, 159, 46, -44),
            (32, 160, 45, -45),
            (33, 161, 44, -46),
            (34, 162, 42, -47),
            (35, 163, 41, -48),
            (36, 164, 40, -49),
            (37, 165, 39, -50),
            (38, 166, 38, -51),
            (39, 167, 36, -52),
            (40, 168, 35, -53),
            (41, 169, 34, -54),
            (42, 170, 32, -55),
            (43, 171, 31, -56),
            (44, 172, 30, -56),
            (45, 173, 28, -57),
            (46, 174, 27, -58),
            (47, 175, 25, -59),
            (48, 176, 24, -59),
            (49, 177, 23, -60),
            (50, 178, 21, -60),
            (51, 179, 20, -61),
            (52, 180, 18, -61),
            (53, 181, 17, -62),
            (54, 182, 15, -62),
            (55, 183, 14, -62),
            (56, 184, 12, -63),
            (57, 185, 10, -63),
            (58, 186, 9, -63),
            (59, 187, 7, -64),
            (60, 188, 6, -64),
            (61, 189, 4, -64),
            (62, 190, 3, -64),
            (63, 191, 1, -64),
            (64, 192, 0, -64),
            (65, 193, -2, -64),
            (66, 194, -3, -64),
            (67, 195, -5, -64),
            (68, 196, -6, -64),
            (69, 197, -8, -64),
            (70, 198, -9, -63),
            (71, 199, -11, -63),
            (72, 200, -12, -63),
            (73, 201, -14, -62),
            (74, 202, -16, -62),
            (75, 203, -17, -62),
            (76, 204, -19, -61),
            (77, 205, -20, -61),
            (78, 206, -22, -60),
            (79, 207, -23, -60),
            (80, 208, -24, -59),
            (81, 209, -26, -59),
            (82, 210, -27, -58),
            (83, 211, -29, -57),
            (84, 212, -30, -56),
            (85, 213, -32, -56),
            (86, 214, -33, -55),
            (87, 215, -34, -54),
            (88, 216, -36, -53),
            (89, 217, -37, -52),
            (90, 218, -38, -51),
            (91, 219, -39, -50),
            (92, 220, -41, -49),
            (93, 221, -42, -48),
            (94, 222, -43, -47),
            (95, 223, -44, -46),
            (96, 224, -45, -45),
            (97, 225, -46, -44),
            (98, 226, -47, -43),
            (99, 227, -48, -42),
            (100, 228, -49, -41),
            (101, 229, -50, -39),
            (102, 230, -51, -38),
            (103, 231, -52, -37),
            (104, 232, -53, -36),
            (105, 233, -54, -34),
            (106, 234, -55, -33),
            (107, 235, -56, -32),
            (108, 236, -56, -30),
            (109, 237, -57, -29),
            (110, 238, -58, -27),
            (111, 239, -59, -26),
            (112, 240, -59, -24),
            (113, 241, -60, -23),
            (114, 242, -60, -22),
            (115, 243, -61, -20),
            (116, 244, -61, -19),
            (117, 245, -62, -17),
            (118, 246, -62, -16),
            (119, 247, -62, -14),
            (120, 248, -63, -12),
            (121, 249, -63, -11),
            (122, 250, -63, -9),
            (123, 251, -64, -8),
            (124, 252, -64, -6),
            (125, 253, -64, -5),
            (126, 254, -64, -3),
            (127, 255, -64, -2));

       signal reg_file : t_data_array(15 downto 0) := (others => (others => '0'));
       signal load_cycles : integer := 0;
       signal run_cycles : integer := 0;
       signal cnt_load : std_logic := '0';
       signal cnt_run  : std_logic := '0';
begin
    
    clock: process
    begin
        clk <= '0';
        clk2x <= '1';
        wait for 5 ns;
        clk2x <= '0';
        wait for 5 ns;
        clk <= '1';
        clk2x <= '1';
        wait for 5 ns;
        clk2x <= '0';
        wait for 5 ns;
    end process clock;

    cnt: process(clk)
    begin
        if rising_edge(clk) then
            if cnt_load = '1' then
                load_cycles <= load_cycles + 1;
            end if;
            if cnt_run = '1' then
                run_cycles <= run_cycles + 1;
            end if;
        end if;
    end process cnt;

    process(clk)
    begin
        if rising_edge(clk) then
            if rst = '0' then
                if reg_ena = '1' then
                    reg_doa <= reg_file(to_integer(unsigned(reg_addra)));
                end if;
                if reg_enb = '1' then
                    reg_dob <= reg_file(to_integer(unsigned(reg_addrb)));
                end if;
            end if;
        end if;
    end process;

    process
        variable l : line;
    begin
        wait for 10 ns;
        wait for 1 ps;
        wait for 40 ns;
        rst <= '0';

        wait for 40 ns;

        prog_cmd(
            (
            arg_type => (
                0 => ARG_IMM,
                1 => ARG_IMM,
                2 => ARG_IMM,
                3 => ARG_IMM,
                4 => ARG_NONE,
                5 => ARG_NONE
            ),
            arg_memchunk => (others => (others => '0')),
            arg_val => (others => '1'),
            arg_assign => (
                0 => "000", -- r
                1 => "001", -- i
                2 => "010", -- addr r
                3 => "011", -- addr i
                4 => "100",
                5 => "101"
            ),
            mem_fetch => (
                0 => '0',
                1 => '0',
                2 => '0',
                3 => '0',
                4 => '0',
                5 => '0'),
            mem_memchunk => (
                0 => "00",
                1 => "00",
                2 => "00",
                3 => "00",
                4 => "00",
                5 => "00"
            ),
            s1_in1a => "000",
            s1_in1b => "000",
            s1_op1  => CALU_NOOP,
            s1_point1 => "000",
            s1_out1 => "000",
            s1_in2a => "000",
            s1_in2b => "000",
            s1_op2 => CALU_NOOP,
            s1_point2 => "000",
            s1_out2 => "000",

            s2_in1a => "000",
            s2_in1b => "000",
            s2_op1  => SALU_NOOP,
            s2_out1 => "000",
            s2_in2a => "000",
            s2_in2b => "000",
            s2_op2  => SALU_NOOP,
            s2_out2  => "000",

            s3_in1a => "000",
            s3_in1b => "000",
            s3_op1  => SALU_NOOP,
            s3_out1 => "000",
            s3_in2a => "000",
            s3_in2b => "000",
            s3_op2  => SALU_NOOP,
            s3_out2 => "000",

            wb => (
                0 => '1',
                1 => '1',
                2 => '0',
                3 => '0',
                4 => '0',
                5 => '0'),
            wb_memchunk => (
                0 => "10", -- R
                1 => "10", -- I
                2 => "00",
                3 => "00",
                4 => "00",
                5 => "00"),
            wb_bitrev => (
                0 => "111",
                1 => "111",
                others => (others => '0')),
            wb_assign => (
                0 => "010",
                1 => "011",
                2 => "000",
                3 => "000",
                4 => "000",
                5 => "000"),
            noop => '0'
            ),
            0,
            start,
            pdata);

        prog_cmd(
            (
            arg_type => (
                0 => ARG_REG, -- i
                1 => ARG_REG, -- j
                2 => ARG_REG, -- r_lut
                3 => ARG_REG, -- i_lut
                4 => ARG_NONE,
                5 => ARG_NONE
            ),
            arg_memchunk => (others => (others => '0')),
            arg_val => (
                0 => '0',
                1 => '0',
                2 => '0',
                3 => '1', -- r_lut
                4 => '1',  -- i_lut
                5 => '0'),
            arg_assign => (
                0 => "000", -- i
                1 => "001", -- j
                2 => "001", -- j
                3 => "010", -- r_lut
                4 => "011", -- i_lut
                5 => "101"),
            mem_fetch => (
                0 => '1',
                1 => '1',
                2 => '1',
                3 => '0',
                4 => '0',
                5 => '0'),
            mem_memchunk => (
                0 => "10", -- R
                1 => "10", -- R
                2 => "11", -- I
                3 => "00",
                4 => "00",
                5 => "00"
            ),
            s1_in1a => "011", -- r_lut
            s1_in1b => "001", -- R[j]
            s1_op1  => CALU_SMUL,
            s1_point1 => "111",
            s1_out1 => "001",
            s1_in2a => "100", -- i_lut
            s1_in2b => "010", -- I[j]
            s1_op2 => CALU_SMUL,
            s1_point2 => "111",
            s1_out2 => "010",

            s2_in1a => "001",
            s2_in1b => "010",
            s2_op1  => SALU_SUB,
            s2_out1 => "001", -- tr
            s2_in2a => "000", -- R[i]
            s2_in2b => ALUIN_1, -- 1
            s2_op2  => SALU_SAR,
            s2_out2  => "000",

            s3_in1a => "000",
            s3_in1b => "001",
            s3_op1  => SALU_SUB,
            s3_out1 => "001",
            s3_in2a => "000",
            s3_in2b => "001",
            s3_op2  => SALU_ADD,
            s3_out2 => "000",

            wb => (
                0 => '1',
                1 => '1',
                2 => '0',
                3 => '0',
                4 => '0',
                5 => '0'),
            wb_memchunk => (
                0 => "10", -- R
                1 => "10", -- R
                2 => "00",
                3 => "00",
                4 => "00",
                5 => "00"),
            wb_bitrev => (others => (others => '0')),
            wb_assign => (
                0 => "000",
                1 => "001",
                2 => "010",
                3 => "011",
                4 => "100",
                5 => "101"),
            noop => '0'
            ),
            1,
            start,
            pdata);

        prog_cmd(
            (
            arg_type => (
                0 => ARG_NONE,
                1 => ARG_NONE,
                2 => ARG_NONE,
                3 => ARG_NONE,
                4 => ARG_NONE,
                5 => ARG_NONE
            ),
            arg_memchunk => (others => (others => '0')),
            arg_val => (others => '0'),
            arg_assign => (
                0 => "000", -- i
                1 => "001", -- j
                2 => "001", -- j
                3 => "010", -- r_lut
                4 => "011", -- i_lut
                5 => "101"
            ),
            mem_fetch => (
                0 => '1',
                1 => '1',
                2 => '1',
                3 => '0',
                4 => '0',
                5 => '0'),
            mem_memchunk => (
                0 => "11", -- I
                1 => "10", -- R
                2 => "11", -- I
                3 => "00",
                4 => "00",
                5 => "00"
            ),
            s1_in1a => "011", -- r_lut
            s1_in1b => "010", -- I[j]
            s1_op1  => CALU_SMUL,
            s1_point1 => "111",
            s1_out1 => "001",
            s1_in2a => "100", -- i_lut
            s1_in2b => "001", -- R[j]
            s1_op2 => CALU_SMUL,
            s1_point2 => "111",
            s1_out2 => "010",

            s2_in1a => "001",
            s2_in1b => "010",
            s2_op1  => SALU_ADD,
            s2_out1 => "001", -- ti
            s2_in2a => "000", -- I[i]
            s2_in2b => ALUIN_1, -- 1
            s2_op2  => SALU_SAR,
            s2_out2  => "000",

            s3_in1a => "000",
            s3_in1b => "001",
            s3_op1  => SALU_SUB,
            s3_out1 => "001",
            s3_in2a => "000",
            s3_in2b => "001",
            s3_op2  => SALU_ADD,
            s3_out2 => "000",

            wb => (
                0 => '1',
                1 => '1',
                2 => '0',
                3 => '0',
                4 => '0',
                5 => '0'),
            wb_memchunk => (
                0 => "11", -- I
                1 => "11", -- I
                2 => "00",
                3 => "00",
                4 => "00",
                5 => "00"),
            wb_bitrev => (others => (others => '0')),
            wb_assign => (
                0 => "000",
                1 => "001",
                2 => "010",
                3 => "011",
                4 => "100",
                5 => "101"),
            noop => '0'
            ),
            2,
            start,
            pdata);

        cnt_load <= '1';
        for i in 0 to 127 loop
            pdata <= "1111111111100000";
            start <= '1';
            wait for 20 ns;
            start <= '0';
            pdata(7 downto 0) <= std_logic_vector(to_signed(sine_wave(i*2), 8));
            pdata(15 downto 8) <= std_logic_vector(to_signed(sine_wave(i*2+1), 8));
            wait for 20 ns;
            pdata(7 downto 0) <= std_logic_vector(to_signed(i*2, 8));
            pdata(15 downto 8) <= std_logic_vector(to_signed(i*2+1, 8));
            wait for 40 ns;
        end loop;
        cnt_load <= '0';

        cnt_run <= '1';
        for i in 0 to 1023 loop
            pdata <= "1111111111100001";
            start <= '1';
            reg_file(0) <= std_logic_vector(to_unsigned(bflys(i)(0), 8));
            reg_file(1) <= std_logic_vector(to_unsigned(bflys(i)(1), 8));
            reg_file(2) <= std_logic_vector(to_signed(bflys(i)(2), 8));
            reg_file(3) <= std_logic_vector(to_signed(bflys(i)(3), 8));
            wait for 20 ns;
            start <= '0';
            pdata(7 downto 0) <= "00000000";
            pdata(15 downto 8) <= "00000001";
            wait for 20 ns;
            pdata(7 downto 0) <= "00000010";
            pdata(15 downto 8) <= "00000011";
            wait for 200 ns;
            pdata <= "1111111111100010";
            start <= '1';
            wait for 20 ns;
            start <= '0';
            wait for 20 ns;
        end loop;
        cnt_run <= '0';

        wait for 140 ns;
        
        mem_ena <= '1';
        mem_enb <= '1';
        for i in 0 to 255 loop
            mem_addra <= "10" & std_logic_vector(to_unsigned(i, 8));
            mem_addrb <= "11" & std_logic_vector(to_unsigned(i, 8));
            wait for 20 ns;
            assert false report integer'image(to_integer(signed(mem_doa))) & ", " & integer'image(to_integer(signed(mem_dob))) severity note;
        end loop;
        mem_ena <= '0';
        mem_enb <= '0';

        wait for 60 ns;

        assert false report "stop load: " & integer'image(load_cycles) & " run: " & integer'image(run_cycles) severity failure;
    end process;
    
    mp_i: entity work.mp
    port map(
        rst => rst,
        clk => clk,
        clk2x => clk2x,
        pdata => pdata,
        pdata_rd => pdata_rd,
        start => start,
        busy => busy,
        mem_addra => mem_addra,
        mem_ena => mem_ena,
        mem_doa => mem_doa,
        mem_addrb => mem_addrb,
        mem_enb => mem_enb,
        mem_dob => mem_dob,
        reg_addra => reg_addra,
        reg_ena => reg_ena,
        reg_doa => reg_doa,
        reg_addrb => reg_addrb,
        reg_enb => reg_enb,
        reg_dob => reg_dob
    );

end behav;
